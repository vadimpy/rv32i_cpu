module top(
    input wire clk,
);



endmodule